module cyberplayer (LSFRout, )